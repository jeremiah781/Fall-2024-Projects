// test.v
module test;
    initial begin
        $display("Icarus Verilog is installed correctly!");
        $finish;
    end
endmodule
