// Testbench for Four-Bit Comparator
//Author: Jeremiah Ddumba
// Date: 2025-01-30
// Description: Simulates the Four-Bit Comparator module with various input combinations.

`timescale 1ns / 1ps

module tb_four_bit_comparator;

// Inputs
reg [3:0] a;
reg [3:0] b;

// Outputs
wire a_equals_b;
wire a_less_than_b;
wire a_greater_than_b;

// Instantiate the Four-Bit Comparator
four_bit_comparator uut (
    .a(a),
    .b(b),
    .a_equals_b(a_equals_b),
    .a_less_than_b(a_less_than_b),
    .a_greater_than_b(a_greater_than_b)
);

integer i, j;

initial begin
    // Display header
    $display("a3 a2 a1 a0 | b3 b2 b1 b0 | eq | lt | gt");
    $display("-------------------------------------------------");
    
    // Iterate through all possible combinations (0 to 15)
    for (i = 0; i < 16; i = i + 1) begin
        for (j = 0; j < 16; j = j + 1) begin
            a = i;
            b = j;
            #1; // Wait for combinational logic to settle
            $display("%b  %b  %b  %b | %b  %b  %b  %b | %b  | %b  | %b",
                     a[3], a[2], a[1], a[0],
                     b[3], b[2], b[1], b[0],
                     a_equals_b, a_less_than_b, a_greater_than_b);
        end
    end
    
    $stop; // End simulation
end

endmodule